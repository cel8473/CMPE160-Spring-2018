library ieee;
use ieee.std_logic_1164.all;

entity T_FF is
port(T, reset, clk : in std_logic;
     Q, QN : inout std_logic := '0');
end T_FF;

architecture behv of T_FF is
begin 
process(reset, clk)
begin
	if(rising_edge(clk)) and reset = '0' then
		if T = '0' then
			Q <= Q after 5 ns;
			QN <= NOT Q after 5 ns; 
		elsif T = '1' then
			Q <= NOT Q after 5 ns;
			QN <= Q after 5 ns;
	elsif reset = '1' then
		Q <= '0' after 5 ns;
		QN <= '1' after 5 ns;
	end if;
	end if;
end process;
end;
