library ieee;
use ieee.std_logic_1164.all;

entity not1 is
port(A : in std_logic;
     Y : out std_logic);
end not1;

architecture df of not1 is
begin
	Y <= NOT A after 4 ns;
end;
