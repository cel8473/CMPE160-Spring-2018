library ieee;
use ieee.std_logic_1164.all;

entity xor3 is
    port(A,B,C : in std_logic;
         Y : out std_logic);
end xor3;

architecture df of xor3 is
begin
  
  Y <= A xor B xor C after 4 ns;
end;

library ieee;
use ieee.std_logic_1164.all;

entity and2 is
  port(A, B : in std_logic;
        Y: out std_logic);
end and2;

architecture df of and2 is 
begin  
  Y <= A AND B after 2 ns;
end;

library ieee;
use ieee.std_logic_1164.all;

entity or3 is 
  port(A, B, C : in std_logic;
       Y: out std_logic);
end or3;

architecture df of or3 is
begin
  Y <= A OR B OR C after 3 ns;
end;